--
--
--  This file is a part of JOP, the Java Optimized Processor
--
--  Copyright (C) 2001-2009, Martin Schoeberl (martin@jopdesign.com)
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--


--
--	microcode.vhd
--
--	Show microcode mnemonic in the simulation
--
--	Author: Peter Hilber
--
--
--
--	2009-08-18	creation
--	FIXME: adapt to new microcode (generate from Instruction.java)
--


library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity microcode is

port (instr : in std_logic_vector(9 downto 0));
end microcode;

architecture sim of microcode is

	type ucval is (
		pop,
		and_uc,
		or_uc,
		xor_uc,
		add,
		sub,
		stmul,
		stmwa,
		stmra,
		stmwd,
		stald,
		stast,
		stgf,
		stpf,
		stcp,
		stbcrd,
		st0,
		st1,
		st2,
		st3,
		st,
		stmi,
		invalid_22,
		invalid_23,
		stvp,
		stjpc,
		star,
		stsp,
		ushr,
		shl,
		shr,
		invalid_31,
		stm_0,
		stm_1,
		stm_2,
		stm_3,
		stm_4,
		stm_5,
		stm_6,
		stm_7,
		stm_8,
		stm_9,
		stm_10,
		stm_11,
		stm_12,
		stm_13,
		stm_14,
		stm_15,
		stm_16,
		stm_17,
		stm_18,
		stm_19,
		stm_20,
		stm_21,
		stm_22,
		stm_23,
		stm_24,
		stm_25,
		stm_26,
		stm_27,
		stm_28,
		stm_29,
		stm_30,
		stm_31,
		bz_idx_0,
		bz_idx_1,
		bz_idx_2,
		bz_idx_3,
		bz_idx_4,
		bz_idx_5,
		bz_idx_6,
		bz_idx_7,
		bz_idx_8,
		bz_idx_9,
		bz_idx_10,
		bz_idx_11,
		bz_idx_12,
		bz_idx_13,
		bz_idx_14,
		bz_idx_15,
		bz_idx_16,
		bz_idx_17,
		bz_idx_18,
		bz_idx_19,
		bz_idx_20,
		bz_idx_21,
		bz_idx_22,
		bz_idx_23,
		bz_idx_24,
		bz_idx_25,
		bz_idx_26,
		bz_idx_27,
		bz_idx_28,
		bz_idx_29,
		bz_idx_30,
		bz_idx_31,
		bnz_idx_0,
		bnz_idx_1,
		bnz_idx_2,
		bnz_idx_3,
		bnz_idx_4,
		bnz_idx_5,
		bnz_idx_6,
		bnz_idx_7,
		bnz_idx_8,
		bnz_idx_9,
		bnz_idx_10,
		bnz_idx_11,
		bnz_idx_12,
		bnz_idx_13,
		bnz_idx_14,
		bnz_idx_15,
		bnz_idx_16,
		bnz_idx_17,
		bnz_idx_18,
		bnz_idx_19,
		bnz_idx_20,
		bnz_idx_21,
		bnz_idx_22,
		bnz_idx_23,
		bnz_idx_24,
		bnz_idx_25,
		bnz_idx_26,
		bnz_idx_27,
		bnz_idx_28,
		bnz_idx_29,
		bnz_idx_30,
		bnz_idx_31,
		nop,
		wait_uc,
		jbr,
		invalid_131,
		invalid_132,
		invalid_133,
		invalid_134,
		invalid_135,
		invalid_136,
		invalid_137,
		invalid_138,
		invalid_139,
		invalid_140,
		invalid_141,
		invalid_142,
		invalid_143,
		invalid_144,
		invalid_145,
		invalid_146,
		invalid_147,
		invalid_148,
		invalid_149,
		invalid_150,
		invalid_151,
		invalid_152,
		invalid_153,
		invalid_154,
		invalid_155,
		invalid_156,
		invalid_157,
		invalid_158,
		invalid_159,
		ldm_0,
		ldm_1,
		ldm_2,
		ldm_3,
		ldm_4,
		ldm_5,
		ldm_6,
		ldm_7,
		ldm_8,
		ldm_9,
		ldm_10,
		ldm_11,
		ldm_12,
		ldm_13,
		ldm_14,
		ldm_15,
		ldm_16,
		ldm_17,
		ldm_18,
		ldm_19,
		ldm_20,
		ldm_21,
		ldm_22,
		ldm_23,
		ldm_24,
		ldm_25,
		ldm_26,
		ldm_27,
		ldm_28,
		ldm_29,
		ldm_30,
		ldm_31,
		ldi_0,
		ldi_1,
		ldi_2,
		ldi_3,
		ldi_4,
		ldi_5,
		ldi_6,
		ldi_7,
		ldi_8,
		ldi_9,
		ldi_10,
		ldi_11,
		ldi_12,
		ldi_13,
		ldi_14,
		ldi_15,
		ldi_16,
		ldi_17,
		ldi_18,
		ldi_19,
		ldi_20,
		ldi_21,
		ldi_22,
		ldi_23,
		ldi_24,
		ldi_25,
		ldi_26,
		ldi_27,
		ldi_28,
		ldi_29,
		ldi_30,
		ldi_31,
		invalid_224,
		invalid_225,
		ldmrd,
		invalid_227,
		invalid_228,
		ldmul,
		invalid_230,
		ldbcstart,
		ld0,
		ld1,
		ld2,
		ld3,
		ld,
		ldmi,
		invalid_238,
		invalid_239,
		ldsp,
		ldvp,
		ldjpc,
		invalid_243,
		ld_opd_8u,
		ld_opd_8s,
		ld_opd_16u,
		ld_opd_16s,
		dup,
		invalid_249,
		invalid_250,
		invalid_251,
		invalid_252,
		invalid_253,
		invalid_254,
		invalid_255			 
	);
	signal val : ucval;

begin

	val <= ucval'val(to_integer(unsigned(instr(7 downto 0))));

end sim;
