--
--
--  This file is a part of JOP, the Java Optimized Processor
--
--  Copyright (C) 2001-2009, Martin Schoeberl (martin@jopdesign.com)
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--


--
--	microcode.vhd
--
--	Show microcode mnemonic in the simulation
--	GENERATED FILE.
--


library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity microcode is

port (instr : in std_logic_vector(9 downto 0));
end microcode;

architecture sim of microcode is

	type ucval is (
		pop,
		and_uc,
		or_uc,
		xor_uc,
		add,
		sub,
		illegal6,
		illegal7,
		illegal8,
		illegal9,
		illegal10,
		illegal11,
		illegal12,
		illegal13,
		illegal14,
		illegal15,
		st0,
		st1,
		st2,
		st3,
		st,
		stmi,
		illegal22,
		illegal23,
		stvp,
		stjpc,
		star,
		stsp,
		ushr,
		shl,
		shr,
		illegal31,
		stm0,
		stm1,
		stm2,
		stm3,
		stm4,
		stm5,
		stm6,
		stm7,
		stm8,
		stm9,
		stm10,
		stm11,
		stm12,
		stm13,
		stm14,
		stm15,
		stm16,
		stm17,
		stm18,
		stm19,
		stm20,
		stm21,
		stm22,
		stm23,
		stm24,
		stm25,
		stm26,
		stm27,
		stm28,
		stm29,
		stm30,
		stm31,
		stmul,
		stmwa,
		stmra,
		stmwd,
		stald,
		stast,
		stgf,
		stpf,
		stcp,
		stbcrd,
		illegal74,
		illegal75,
		illegal76,
		illegal77,
		illegal78,
		illegal79,
		illegal80,
		illegal81,
		illegal82,
		illegal83,
		illegal84,
		illegal85,
		illegal86,
		illegal87,
		illegal88,
		illegal89,
		illegal90,
		illegal91,
		illegal92,
		illegal93,
		illegal94,
		illegal95,
		illegal96,
		illegal97,
		illegal98,
		illegal99,
		illegal100,
		illegal101,
		illegal102,
		illegal103,
		illegal104,
		illegal105,
		illegal106,
		illegal107,
		illegal108,
		illegal109,
		illegal110,
		illegal111,
		illegal112,
		illegal113,
		illegal114,
		illegal115,
		illegal116,
		illegal117,
		illegal118,
		illegal119,
		illegal120,
		illegal121,
		illegal122,
		illegal123,
		illegal124,
		illegal125,
		illegal126,
		illegal127,
		illegal128,
		illegal129,
		illegal130,
		illegal131,
		illegal132,
		illegal133,
		illegal134,
		illegal135,
		illegal136,
		illegal137,
		illegal138,
		illegal139,
		illegal140,
		illegal141,
		illegal142,
		illegal143,
		illegal144,
		illegal145,
		illegal146,
		illegal147,
		illegal148,
		illegal149,
		illegal150,
		illegal151,
		illegal152,
		illegal153,
		illegal154,
		illegal155,
		illegal156,
		illegal157,
		illegal158,
		illegal159,
		ldm0,
		ldm1,
		ldm2,
		ldm3,
		ldm4,
		ldm5,
		ldm6,
		ldm7,
		ldm8,
		ldm9,
		ldm10,
		ldm11,
		ldm12,
		ldm13,
		ldm14,
		ldm15,
		ldm16,
		ldm17,
		ldm18,
		ldm19,
		ldm20,
		ldm21,
		ldm22,
		ldm23,
		ldm24,
		ldm25,
		ldm26,
		ldm27,
		ldm28,
		ldm29,
		ldm30,
		ldm31,
		ldi0,
		ldi1,
		ldi2,
		ldi3,
		ldi4,
		ldi5,
		ldi6,
		ldi7,
		ldi8,
		ldi9,
		ldi10,
		ldi11,
		ldi12,
		ldi13,
		ldi14,
		ldi15,
		ldi16,
		ldi17,
		ldi18,
		ldi19,
		ldi20,
		ldi21,
		ldi22,
		ldi23,
		ldi24,
		ldi25,
		ldi26,
		ldi27,
		ldi28,
		ldi29,
		ldi30,
		ldi31,
		ldmrd,
		ldmul,
		ldbcstart,
		illegal227,
		illegal228,
		illegal229,
		illegal230,
		illegal231,
		ld0,
		ld1,
		ld2,
		ld3,
		ld,
		ldmi,
		illegal238,
		illegal239,
		ldsp,
		ldvp,
		ldjpc,
		illegal243,
		ld_opd_8u,
		ld_opd_8s,
		ld_opd_16u,
		ld_opd_16s,
		dup,
		illegal249,
		illegal250,
		illegal251,
		illegal252,
		illegal253,
		illegal254,
		illegal255,
		nop,
		wait_uc,
		jbr,
		illegal259,
		illegal260,
		illegal261,
		illegal262,
		illegal263,
		illegal264,
		illegal265,
		illegal266,
		illegal267,
		illegal268,
		illegal269,
		illegal270,
		illegal271,
		illegal272,
		illegal273,
		illegal274,
		illegal275,
		illegal276,
		illegal277,
		illegal278,
		illegal279,
		illegal280,
		illegal281,
		illegal282,
		illegal283,
		illegal284,
		illegal285,
		illegal286,
		illegal287,
		illegal288,
		illegal289,
		illegal290,
		illegal291,
		illegal292,
		illegal293,
		illegal294,
		illegal295,
		illegal296,
		illegal297,
		illegal298,
		illegal299,
		illegal300,
		illegal301,
		illegal302,
		illegal303,
		illegal304,
		illegal305,
		illegal306,
		illegal307,
		illegal308,
		illegal309,
		illegal310,
		illegal311,
		illegal312,
		illegal313,
		illegal314,
		illegal315,
		illegal316,
		illegal317,
		illegal318,
		illegal319,
		illegal320,
		illegal321,
		illegal322,
		illegal323,
		illegal324,
		illegal325,
		illegal326,
		illegal327,
		illegal328,
		illegal329,
		illegal330,
		illegal331,
		illegal332,
		illegal333,
		illegal334,
		illegal335,
		illegal336,
		illegal337,
		illegal338,
		illegal339,
		illegal340,
		illegal341,
		illegal342,
		illegal343,
		illegal344,
		illegal345,
		illegal346,
		illegal347,
		illegal348,
		illegal349,
		illegal350,
		illegal351,
		illegal352,
		illegal353,
		illegal354,
		illegal355,
		illegal356,
		illegal357,
		illegal358,
		illegal359,
		illegal360,
		illegal361,
		illegal362,
		illegal363,
		illegal364,
		illegal365,
		illegal366,
		illegal367,
		illegal368,
		illegal369,
		illegal370,
		illegal371,
		illegal372,
		illegal373,
		illegal374,
		illegal375,
		illegal376,
		illegal377,
		illegal378,
		illegal379,
		illegal380,
		illegal381,
		illegal382,
		illegal383,
		bz0,
		bz1,
		bz2,
		bz3,
		bz4,
		bz5,
		bz6,
		bz7,
		bz8,
		bz9,
		bz10,
		bz11,
		bz12,
		bz13,
		bz14,
		bz15,
		bz16,
		bz17,
		bz18,
		bz19,
		bz20,
		bz21,
		bz22,
		bz23,
		bz24,
		bz25,
		bz26,
		bz27,
		bz28,
		bz29,
		bz30,
		bz31,
		bz32,
		bz33,
		bz34,
		bz35,
		bz36,
		bz37,
		bz38,
		bz39,
		bz40,
		bz41,
		bz42,
		bz43,
		bz44,
		bz45,
		bz46,
		bz47,
		bz48,
		bz49,
		bz50,
		bz51,
		bz52,
		bz53,
		bz54,
		bz55,
		bz56,
		bz57,
		bz58,
		bz59,
		bz60,
		bz61,
		bz62,
		bz63,
		bnz0,
		bnz1,
		bnz2,
		bnz3,
		bnz4,
		bnz5,
		bnz6,
		bnz7,
		bnz8,
		bnz9,
		bnz10,
		bnz11,
		bnz12,
		bnz13,
		bnz14,
		bnz15,
		bnz16,
		bnz17,
		bnz18,
		bnz19,
		bnz20,
		bnz21,
		bnz22,
		bnz23,
		bnz24,
		bnz25,
		bnz26,
		bnz27,
		bnz28,
		bnz29,
		bnz30,
		bnz31,
		bnz32,
		bnz33,
		bnz34,
		bnz35,
		bnz36,
		bnz37,
		bnz38,
		bnz39,
		bnz40,
		bnz41,
		bnz42,
		bnz43,
		bnz44,
		bnz45,
		bnz46,
		bnz47,
		bnz48,
		bnz49,
		bnz50,
		bnz51,
		bnz52,
		bnz53,
		bnz54,
		bnz55,
		bnz56,
		bnz57,
		bnz58,
		bnz59,
		bnz60,
		bnz61,
		bnz62,
		bnz63,
		jmp0,
		jmp1,
		jmp2,
		jmp3,
		jmp4,
		jmp5,
		jmp6,
		jmp7,
		jmp8,
		jmp9,
		jmp10,
		jmp11,
		jmp12,
		jmp13,
		jmp14,
		jmp15,
		jmp16,
		jmp17,
		jmp18,
		jmp19,
		jmp20,
		jmp21,
		jmp22,
		jmp23,
		jmp24,
		jmp25,
		jmp26,
		jmp27,
		jmp28,
		jmp29,
		jmp30,
		jmp31,
		jmp32,
		jmp33,
		jmp34,
		jmp35,
		jmp36,
		jmp37,
		jmp38,
		jmp39,
		jmp40,
		jmp41,
		jmp42,
		jmp43,
		jmp44,
		jmp45,
		jmp46,
		jmp47,
		jmp48,
		jmp49,
		jmp50,
		jmp51,
		jmp52,
		jmp53,
		jmp54,
		jmp55,
		jmp56,
		jmp57,
		jmp58,
		jmp59,
		jmp60,
		jmp61,
		jmp62,
		jmp63,
		jmp64,
		jmp65,
		jmp66,
		jmp67,
		jmp68,
		jmp69,
		jmp70,
		jmp71,
		jmp72,
		jmp73,
		jmp74,
		jmp75,
		jmp76,
		jmp77,
		jmp78,
		jmp79,
		jmp80,
		jmp81,
		jmp82,
		jmp83,
		jmp84,
		jmp85,
		jmp86,
		jmp87,
		jmp88,
		jmp89,
		jmp90,
		jmp91,
		jmp92,
		jmp93,
		jmp94,
		jmp95,
		jmp96,
		jmp97,
		jmp98,
		jmp99,
		jmp100,
		jmp101,
		jmp102,
		jmp103,
		jmp104,
		jmp105,
		jmp106,
		jmp107,
		jmp108,
		jmp109,
		jmp110,
		jmp111,
		jmp112,
		jmp113,
		jmp114,
		jmp115,
		jmp116,
		jmp117,
		jmp118,
		jmp119,
		jmp120,
		jmp121,
		jmp122,
		jmp123,
		jmp124,
		jmp125,
		jmp126,
		jmp127,
		jmp128,
		jmp129,
		jmp130,
		jmp131,
		jmp132,
		jmp133,
		jmp134,
		jmp135,
		jmp136,
		jmp137,
		jmp138,
		jmp139,
		jmp140,
		jmp141,
		jmp142,
		jmp143,
		jmp144,
		jmp145,
		jmp146,
		jmp147,
		jmp148,
		jmp149,
		jmp150,
		jmp151,
		jmp152,
		jmp153,
		jmp154,
		jmp155,
		jmp156,
		jmp157,
		jmp158,
		jmp159,
		jmp160,
		jmp161,
		jmp162,
		jmp163,
		jmp164,
		jmp165,
		jmp166,
		jmp167,
		jmp168,
		jmp169,
		jmp170,
		jmp171,
		jmp172,
		jmp173,
		jmp174,
		jmp175,
		jmp176,
		jmp177,
		jmp178,
		jmp179,
		jmp180,
		jmp181,
		jmp182,
		jmp183,
		jmp184,
		jmp185,
		jmp186,
		jmp187,
		jmp188,
		jmp189,
		jmp190,
		jmp191,
		jmp192,
		jmp193,
		jmp194,
		jmp195,
		jmp196,
		jmp197,
		jmp198,
		jmp199,
		jmp200,
		jmp201,
		jmp202,
		jmp203,
		jmp204,
		jmp205,
		jmp206,
		jmp207,
		jmp208,
		jmp209,
		jmp210,
		jmp211,
		jmp212,
		jmp213,
		jmp214,
		jmp215,
		jmp216,
		jmp217,
		jmp218,
		jmp219,
		jmp220,
		jmp221,
		jmp222,
		jmp223,
		jmp224,
		jmp225,
		jmp226,
		jmp227,
		jmp228,
		jmp229,
		jmp230,
		jmp231,
		jmp232,
		jmp233,
		jmp234,
		jmp235,
		jmp236,
		jmp237,
		jmp238,
		jmp239,
		jmp240,
		jmp241,
		jmp242,
		jmp243,
		jmp244,
		jmp245,
		jmp246,
		jmp247,
		jmp248,
		jmp249,
		jmp250,
		jmp251,
		jmp252,
		jmp253,
		jmp254,
		jmp255,
		jmp256,
		jmp257,
		jmp258,
		jmp259,
		jmp260,
		jmp261,
		jmp262,
		jmp263,
		jmp264,
		jmp265,
		jmp266,
		jmp267,
		jmp268,
		jmp269,
		jmp270,
		jmp271,
		jmp272,
		jmp273,
		jmp274,
		jmp275,
		jmp276,
		jmp277,
		jmp278,
		jmp279,
		jmp280,
		jmp281,
		jmp282,
		jmp283,
		jmp284,
		jmp285,
		jmp286,
		jmp287,
		jmp288,
		jmp289,
		jmp290,
		jmp291,
		jmp292,
		jmp293,
		jmp294,
		jmp295,
		jmp296,
		jmp297,
		jmp298,
		jmp299,
		jmp300,
		jmp301,
		jmp302,
		jmp303,
		jmp304,
		jmp305,
		jmp306,
		jmp307,
		jmp308,
		jmp309,
		jmp310,
		jmp311,
		jmp312,
		jmp313,
		jmp314,
		jmp315,
		jmp316,
		jmp317,
		jmp318,
		jmp319,
		jmp320,
		jmp321,
		jmp322,
		jmp323,
		jmp324,
		jmp325,
		jmp326,
		jmp327,
		jmp328,
		jmp329,
		jmp330,
		jmp331,
		jmp332,
		jmp333,
		jmp334,
		jmp335,
		jmp336,
		jmp337,
		jmp338,
		jmp339,
		jmp340,
		jmp341,
		jmp342,
		jmp343,
		jmp344,
		jmp345,
		jmp346,
		jmp347,
		jmp348,
		jmp349,
		jmp350,
		jmp351,
		jmp352,
		jmp353,
		jmp354,
		jmp355,
		jmp356,
		jmp357,
		jmp358,
		jmp359,
		jmp360,
		jmp361,
		jmp362,
		jmp363,
		jmp364,
		jmp365,
		jmp366,
		jmp367,
		jmp368,
		jmp369,
		jmp370,
		jmp371,
		jmp372,
		jmp373,
		jmp374,
		jmp375,
		jmp376,
		jmp377,
		jmp378,
		jmp379,
		jmp380,
		jmp381,
		jmp382,
		jmp383,
		jmp384,
		jmp385,
		jmp386,
		jmp387,
		jmp388,
		jmp389,
		jmp390,
		jmp391,
		jmp392,
		jmp393,
		jmp394,
		jmp395,
		jmp396,
		jmp397,
		jmp398,
		jmp399,
		jmp400,
		jmp401,
		jmp402,
		jmp403,
		jmp404,
		jmp405,
		jmp406,
		jmp407,
		jmp408,
		jmp409,
		jmp410,
		jmp411,
		jmp412,
		jmp413,
		jmp414,
		jmp415,
		jmp416,
		jmp417,
		jmp418,
		jmp419,
		jmp420,
		jmp421,
		jmp422,
		jmp423,
		jmp424,
		jmp425,
		jmp426,
		jmp427,
		jmp428,
		jmp429,
		jmp430,
		jmp431,
		jmp432,
		jmp433,
		jmp434,
		jmp435,
		jmp436,
		jmp437,
		jmp438,
		jmp439,
		jmp440,
		jmp441,
		jmp442,
		jmp443,
		jmp444,
		jmp445,
		jmp446,
		jmp447,
		jmp448,
		jmp449,
		jmp450,
		jmp451,
		jmp452,
		jmp453,
		jmp454,
		jmp455,
		jmp456,
		jmp457,
		jmp458,
		jmp459,
		jmp460,
		jmp461,
		jmp462,
		jmp463,
		jmp464,
		jmp465,
		jmp466,
		jmp467,
		jmp468,
		jmp469,
		jmp470,
		jmp471,
		jmp472,
		jmp473,
		jmp474,
		jmp475,
		jmp476,
		jmp477,
		jmp478,
		jmp479,
		jmp480,
		jmp481,
		jmp482,
		jmp483,
		jmp484,
		jmp485,
		jmp486,
		jmp487,
		jmp488,
		jmp489,
		jmp490,
		jmp491,
		jmp492,
		jmp493,
		jmp494,
		jmp495,
		jmp496,
		jmp497,
		jmp498,
		jmp499,
		jmp500,
		jmp501,
		jmp502,
		jmp503,
		jmp504,
		jmp505,
		jmp506,
		jmp507,
		jmp508,
		jmp509,
		jmp510,
		jmp511
);
	signal val : ucval;

begin

	val <= ucval'val(to_integer(unsigned(instr)));

end sim;
