--
--
--  This file is a part of JOP, the Java Optimized Processor
--
--  Copyright (C) 2009, Martin Schoeberl (martin@jopdesign.com)
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--


--
--	microcode.vhd
--
--	Show microcode mnemonic in the simulation
--
--	Author: Peter Hilber, Martin Schoeberl
--
--
--	2009-08-18	creation
--	2009-11-25	generate the mnemonics from Instruction.java
--


library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity microcode is

port (instr : in std_logic_vector(9 downto 0));
end microcode;

architecture sim of microcode is

-- the following code is generated by Instruction.java ---------

	type mcval is (
		pop,
		and_x,
		or_x,
		xor_x,
		add,
		sub,
		st0,
		st1,
		st2,
		st3,
		st,
		stmi,
		stvp,
		stjpc,
		star,
		stsp,
		ushr,
		shl,
		shr,
		stm,
		stmul,
		stmwa,
		stmra,
		stmwd,
		stald,
		stast,
		stgf,
		stpf,
		stcp,
		stbcrd,
		stidx,
		stps,
		stmrac,
		stmraf,
		stmwdf,
		ldm,
		ldi,
		ldmrd,
		ldmul,
		ldbcstart,
		ld0,
		ld1,
		ld2,
		ld3,
		ld,
		ldmi,
		ldsp,
		ldvp,
		ldjpc,
		ld_opd_8u,
		ld_opd_8s,
		ld_opd_16u,
		ld_opd_16s,
		dup,
		nop,
		wait_x,
		jbr,
		stgs,
		bz,
		bnz,
		jmp,
		unknown
	);
	signal val : mcval;


begin

process(instr)
begin

	val <= unknown;
	if instr(9)='1' then
		val <= jmp;
	elsif instr(9 downto 6)="0110" then
		val <= bz;
	elsif instr(9 downto 6)="0111" then
		val <= bnz;
	else
		case instr is
			when "0000000000" => val <= pop;
			when "0000000001" => val <= and_x;
			when "0000000010" => val <= or_x;
			when "0000000011" => val <= xor_x;
			when "0000000100" => val <= add;
			when "0000000101" => val <= sub;
			when "0000010000" => val <= st0;
			when "0000010001" => val <= st1;
			when "0000010010" => val <= st2;
			when "0000010011" => val <= st3;
			when "0000010100" => val <= st;
			when "0000010101" => val <= stmi;
			when "0000011000" => val <= stvp;
			when "0000011001" => val <= stjpc;
			when "0000011010" => val <= star;
			when "0000011011" => val <= stsp;
			when "0000011100" => val <= ushr;
			when "0000011101" => val <= shl;
			when "0000011110" => val <= shr;
			when "0000100000" => val <= stm;
			when "0000100001" => val <= stm;
			when "0000100010" => val <= stm;
			when "0000100011" => val <= stm;
			when "0000100100" => val <= stm;
			when "0000100101" => val <= stm;
			when "0000100110" => val <= stm;
			when "0000100111" => val <= stm;
			when "0000101000" => val <= stm;
			when "0000101001" => val <= stm;
			when "0000101010" => val <= stm;
			when "0000101011" => val <= stm;
			when "0000101100" => val <= stm;
			when "0000101101" => val <= stm;
			when "0000101110" => val <= stm;
			when "0000101111" => val <= stm;
			when "0000110000" => val <= stm;
			when "0000110001" => val <= stm;
			when "0000110010" => val <= stm;
			when "0000110011" => val <= stm;
			when "0000110100" => val <= stm;
			when "0000110101" => val <= stm;
			when "0000110110" => val <= stm;
			when "0000110111" => val <= stm;
			when "0000111000" => val <= stm;
			when "0000111001" => val <= stm;
			when "0000111010" => val <= stm;
			when "0000111011" => val <= stm;
			when "0000111100" => val <= stm;
			when "0000111101" => val <= stm;
			when "0000111110" => val <= stm;
			when "0000111111" => val <= stm;
			when "0001000000" => val <= stmul;
			when "0001000001" => val <= stmwa;
			when "0001000010" => val <= stmra;
			when "0001000011" => val <= stmwd;
			when "0001000100" => val <= stald;
			when "0001000101" => val <= stast;
			when "0001000110" => val <= stgf;
			when "0001000111" => val <= stpf;
			when "0001001000" => val <= stcp;
			when "0001001001" => val <= stbcrd;
			when "0001001010" => val <= stidx;
			when "0001001011" => val <= stps;
			when "0001001100" => val <= stmrac;
			when "0001001101" => val <= stmraf;
			when "0001001110" => val <= stmwdf;
			when "0010100000" => val <= ldm;
			when "0010100001" => val <= ldm;
			when "0010100010" => val <= ldm;
			when "0010100011" => val <= ldm;
			when "0010100100" => val <= ldm;
			when "0010100101" => val <= ldm;
			when "0010100110" => val <= ldm;
			when "0010100111" => val <= ldm;
			when "0010101000" => val <= ldm;
			when "0010101001" => val <= ldm;
			when "0010101010" => val <= ldm;
			when "0010101011" => val <= ldm;
			when "0010101100" => val <= ldm;
			when "0010101101" => val <= ldm;
			when "0010101110" => val <= ldm;
			when "0010101111" => val <= ldm;
			when "0010110000" => val <= ldm;
			when "0010110001" => val <= ldm;
			when "0010110010" => val <= ldm;
			when "0010110011" => val <= ldm;
			when "0010110100" => val <= ldm;
			when "0010110101" => val <= ldm;
			when "0010110110" => val <= ldm;
			when "0010110111" => val <= ldm;
			when "0010111000" => val <= ldm;
			when "0010111001" => val <= ldm;
			when "0010111010" => val <= ldm;
			when "0010111011" => val <= ldm;
			when "0010111100" => val <= ldm;
			when "0010111101" => val <= ldm;
			when "0010111110" => val <= ldm;
			when "0010111111" => val <= ldm;
			when "0011000000" => val <= ldi;
			when "0011000001" => val <= ldi;
			when "0011000010" => val <= ldi;
			when "0011000011" => val <= ldi;
			when "0011000100" => val <= ldi;
			when "0011000101" => val <= ldi;
			when "0011000110" => val <= ldi;
			when "0011000111" => val <= ldi;
			when "0011001000" => val <= ldi;
			when "0011001001" => val <= ldi;
			when "0011001010" => val <= ldi;
			when "0011001011" => val <= ldi;
			when "0011001100" => val <= ldi;
			when "0011001101" => val <= ldi;
			when "0011001110" => val <= ldi;
			when "0011001111" => val <= ldi;
			when "0011010000" => val <= ldi;
			when "0011010001" => val <= ldi;
			when "0011010010" => val <= ldi;
			when "0011010011" => val <= ldi;
			when "0011010100" => val <= ldi;
			when "0011010101" => val <= ldi;
			when "0011010110" => val <= ldi;
			when "0011010111" => val <= ldi;
			when "0011011000" => val <= ldi;
			when "0011011001" => val <= ldi;
			when "0011011010" => val <= ldi;
			when "0011011011" => val <= ldi;
			when "0011011100" => val <= ldi;
			when "0011011101" => val <= ldi;
			when "0011011110" => val <= ldi;
			when "0011011111" => val <= ldi;
			when "0011100000" => val <= ldmrd;
			when "0011100001" => val <= ldmul;
			when "0011100010" => val <= ldbcstart;
			when "0011101000" => val <= ld0;
			when "0011101001" => val <= ld1;
			when "0011101010" => val <= ld2;
			when "0011101011" => val <= ld3;
			when "0011101100" => val <= ld;
			when "0011101101" => val <= ldmi;
			when "0011110000" => val <= ldsp;
			when "0011110001" => val <= ldvp;
			when "0011110010" => val <= ldjpc;
			when "0011110100" => val <= ld_opd_8u;
			when "0011110101" => val <= ld_opd_8s;
			when "0011110110" => val <= ld_opd_16u;
			when "0011110111" => val <= ld_opd_16s;
			when "0011111000" => val <= dup;
			when "0100000000" => val <= nop;
			when "0100000001" => val <= wait_x;
			when "0100000010" => val <= jbr;
			when "0100010000" => val <= stgs;

			when others => null;
		end case;
	end if;

end process;

-- end generated code ------------------------------------------

end sim;
