-- pragma translate_off
use std.textio.all;
-- pragma translate_on
package version is
  constant grlib_version : integer := 1014;
-- pragma translate_off
  constant grlib_date : string := "20070227";
-- pragma translate_on
  constant grlib_build : integer := 2053;
end;
