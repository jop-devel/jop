--
--  This file is part of JOP, the Java Optimized Processor
--
--  Copyright (C) 2007,2008, Christof Pitter
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.sc_pack.all;

package sc_arbiter_pack is
	
	type arb_out_type is array (integer range <>) of sc_out_type;
	type arb_in_type is array (integer range <>) of sc_in_type;
	
	-- TM
	
	type tm_broadcast_type is record
		valid : std_logic;
		address : std_logic_vector(SC_ADDR_SIZE-1 downto 0);
	end record; 

end sc_arbiter_pack;
