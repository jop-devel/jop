pll_inst : pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
