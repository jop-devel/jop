--
--	jop_types_20.vhd
--
--	package for 20MHz definitions
--


package jop_types is

	-- constants for 20MHz input and 20MHz internal clock
	constant clk_freq : integer := 20000000;
	constant pll_mult : natural := 1;
	constant pll_div : natural := 1;

end jop_types;

package body jop_types is

end jop_types;
